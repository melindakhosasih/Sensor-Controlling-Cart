module SevenSegment(
	output reg [6:0] display,
	output reg [3:0] digit,
	input wire [15:0] nums,
	input wire rst,
	input wire clk
    );
    
    reg [15:0] clk_divider;
    reg [3:0] display_num;
    
    always @ (posedge clk) begin
    	clk_divider <= clk_divider + 15'b1;
    end
    
    always @ (posedge clk_divider[15]) begin
		case (digit)
			4'b1110 : begin
					display_num <= nums[7:4];
					digit <= 4'b1101;
				end
			4'b1101 : begin
					display_num <= nums[11:8];
					digit <= 4'b1011;
				end
			4'b1011 : begin
					display_num <= nums[15:12];
					digit <= 4'b0111;
				end
			4'b0111 : begin
					display_num <= nums[3:0];
					digit <= 4'b1110;
				end
			default : begin
					display_num <= nums[3:0];
					digit <= 4'b1110;
				end				
		endcase
    end
    
    always @ (*) begin
    	case (display_num)
    		0 : display = 7'b1000000;	//0000
			1 : display = 7'b1111001;   //0001                                                
			2 : display = 7'b0100100;   //0010                                                
			3 : display = 7'b0110000;   //0011                                             
			4 : display = 7'b0011001;   //0100                                               
			5 : display = 7'b0010010;   //0101                                               
			6 : display = 7'b0000010;   //0110
			7 : display = 7'b1111000;   //0111
			8 : display = 7'b0000000;   //1000
			9 : display = 7'b0010000;	//1001
			default : display = 7'b1111111;
    	endcase
    end
    
endmodule
